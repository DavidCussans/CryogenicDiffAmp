.title KiCad schematic
Rqp1 /cathode /N002 {Rq / Np }
Cqp1 /cathode /N002 {Cq * Np}
Cdp1 /N002 /anode {Cd * Np}
Rq1 /cathode /N001 {Rq / Nf }
Cq1 /cathode /N001 {Cq * Nf}
Cd1 /N001 /anode {Cd * Nf}
Vbd1 /N006 /anode dc 70
Vtr1 /N005 /N006 dc 400m
Rd1 /N006 /N004 {Rd/Nf}
Cg1 /cathode /anode {Cg}
SQuench1 /N001 /N004 /N003 PSpiceSwitch
U1 /N004 /N005 /N003 AMP
STrigger1 /N001 /N004 0 PSpiceSwitch
.SUBCKT SiPMT  /anode /cathode /ph Cd=80f Cq=8f Cm=59p Cg=59p Rd=1k Rq=300k Nf=1 Np=3599 Ith=100u Vbd=70.5
.ends
.end
