.title KiCad schematic
.include "../SiPMT_model2.cir"
V2 Net-_D1-Pad3_ 0 dc 0 ac 0 pulse(0V 1V 10n 1n 1n 1n)
XD1 /va /vk Net-_D1-Pad3_ SiPMT Np=35990
R2 /va 0 50
V1 /vk 0 72.0
.control
option savecurrents
tran 1ns 100ns
write
.endc
.end
